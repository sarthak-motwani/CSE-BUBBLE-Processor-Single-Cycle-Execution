
module InstMem(clock, address, inst);

	input clock;
	input [31:0] address;
	
	output reg [31:0]	inst;
	
	reg [31:0] Mem [0:127];
	
	initial begin
	
		Mem[1] = 32'b00000000001001010010100000100000;
		Mem[0] = 32'b00000000100000000010100000100000;
		Mem[2] = 32'b10001100101001100000000000000000;
		Mem[3] = 32'b10001100101001110000000000000001;
		Mem[4] = 32'b00000000110001110100000000101010;
		Mem[5] = 32'b00010101000000000000000000000010;
		Mem[6] = 32'b10101100101001110000000000000000;
		Mem[7] = 32'b10101100101001100000000000000001;
		Mem[8] = 32'b00100000100001000000000000000001;
		Mem[9] = 32'b00000000011000100100100000100010;
		Mem[10] = 32'b00010100100010011111111111110101;
		Mem[11] = 32'b00100000010000100000000000000001;
		Mem[12] = 32'b10001100000001000000000000000000;
		Mem[13] = 32'b00010100010000111111111111110010;
	

	end
	
	always @( posedge clock) begin
		inst <= Mem[address[6:0]];
	end
endmodule